module prob1d (inA, inB, out);

input [7:0] inA, inB;
output [8:0] out;

assign out = inA + inB;

endmodule